-- embedded_computer_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity embedded_computer_system is
	port (
		buffer_1_call_valid         : in    std_logic                     := '0';             --        buffer_1_call.valid
		buffer_1_call_stall         : out   std_logic;                                        --                     .stall
		buffer_1_return_valid       : out   std_logic;                                        --      buffer_1_return.valid
		buffer_1_return_stall       : in    std_logic                     := '0';             --                     .stall
		clk_clk                     : in    std_logic                     := '0';             --                  clk.clk
		filter_0_call_valid         : in    std_logic                     := '0';             --        filter_0_call.valid
		filter_0_call_stall         : out   std_logic;                                        --                     .stall
		filter_0_return_valid       : out   std_logic;                                        --      filter_0_return.valid
		filter_0_return_stall       : in    std_logic                     := '0';             --                     .stall
		pll_c1_clk                  : out   std_logic;                                        --               pll_c1.clk
		reset_reset_n               : in    std_logic                     := '0';             --                reset.reset_n
		sdram_controller_addr       : out   std_logic_vector(12 downto 0);                    --     sdram_controller.addr
		sdram_controller_ba         : out   std_logic_vector(1 downto 0);                     --                     .ba
		sdram_controller_cas_n      : out   std_logic;                                        --                     .cas_n
		sdram_controller_cke        : out   std_logic;                                        --                     .cke
		sdram_controller_cs_n       : out   std_logic;                                        --                     .cs_n
		sdram_controller_dq         : inout std_logic_vector(15 downto 0) := (others => '0'); --                     .dq
		sdram_controller_dqm        : out   std_logic_vector(1 downto 0);                     --                     .dqm
		sdram_controller_ras_n      : out   std_logic;                                        --                     .ras_n
		sdram_controller_we_n       : out   std_logic;                                        --                     .we_n
		vga_ip_0_conduit_end_vga_b  : out   std_logic_vector(3 downto 0);                     -- vga_ip_0_conduit_end.vga_b
		vga_ip_0_conduit_end_vga_g  : out   std_logic_vector(3 downto 0);                     --                     .vga_g
		vga_ip_0_conduit_end_vga_r  : out   std_logic_vector(3 downto 0);                     --                     .vga_r
		vga_ip_0_conduit_end_vga_vs : out   std_logic;                                        --                     .vga_vs
		vga_ip_0_conduit_end_vga_hs : out   std_logic                                         --                     .vga_hs
	);
end entity embedded_computer_system;

architecture rtl of embedded_computer_system is
	component TIMER_HW_IP is
		port (
			reset_n : in  std_logic                     := 'X';             -- reset_n
			clk     : in  std_logic                     := 'X';             -- clk
			cs_n    : in  std_logic                     := 'X';             -- chipselect_n
			addr    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n : in  std_logic                     := 'X';             -- write_n
			read_n  : in  std_logic                     := 'X';             -- read_n
			din     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dout    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component TIMER_HW_IP;

	component VGA_IP is
		port (
			data_controller_in    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wren_controller       : in  std_logic                     := 'X';             -- write
			cs_n                  : in  std_logic                     := 'X';             -- chipselect_n
			address_controller_in : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			reset_controller      : in  std_logic                     := 'X';             -- reset_n
			CLOCK_controller_50   : in  std_logic                     := 'X';             -- clk
			VGA_controller_B      : out std_logic_vector(3 downto 0);                     -- vga_b
			VGA_controller_G      : out std_logic_vector(3 downto 0);                     -- vga_g
			VGA_controller_R      : out std_logic_vector(3 downto 0);                     -- vga_r
			VGA_controller_VS     : out std_logic;                                        -- vga_vs
			VGA_controller_HS     : out std_logic                                         -- vga_hs
		);
	end component VGA_IP;

	component embedded_computer_system_buffer_0 is
		port (
			avs_cra_read                 : in  std_logic                     := 'X';             -- read
			avs_cra_write                : in  std_logic                     := 'X';             -- write
			avs_cra_address              : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avs_cra_writedata            : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cra_byteenable           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avs_cra_readdata             : out std_logic_vector(63 downto 0);                    -- readdata
			avs_sample_buffer_read       : in  std_logic                     := 'X';             -- read
			avs_sample_buffer_write      : in  std_logic                     := 'X';             -- write
			avs_sample_buffer_address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			avs_sample_buffer_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_sample_buffer_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_sample_buffer_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			clock                        : in  std_logic                     := 'X';             -- clk
			done_irq                     : out std_logic;                                        -- irq
			resetn                       : in  std_logic                     := 'X';             -- reset_n
			sample_out_data              : out std_logic_vector(15 downto 0);                    -- data
			sample_out_ready             : in  std_logic                     := 'X';             -- ready
			sample_out_valid             : out std_logic                                         -- valid
		);
	end component embedded_computer_system_buffer_0;

	component embedded_computer_system_buffer_1 is
		port (
			avs_result_buffer_read       : in  std_logic                     := 'X';             -- read
			avs_result_buffer_write      : in  std_logic                     := 'X';             -- write
			avs_result_buffer_address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			avs_result_buffer_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_result_buffer_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_result_buffer_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			start                        : in  std_logic                     := 'X';             -- valid
			busy                         : out std_logic;                                        -- stall
			clock                        : in  std_logic                     := 'X';             -- clk
			resetn                       : in  std_logic                     := 'X';             -- reset_n
			result_in_data               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			result_in_ready              : out std_logic;                                        -- ready
			result_in_valid              : in  std_logic                     := 'X';             -- valid
			done                         : out std_logic;                                        -- valid
			stall                        : in  std_logic                     := 'X'              -- stall
		);
	end component embedded_computer_system_buffer_1;

	component embedded_computer_system_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component embedded_computer_system_cpu;

	component embedded_computer_system_filter_0 is
		port (
			start         : in  std_logic                     := 'X';             -- valid
			busy          : out std_logic;                                        -- stall
			clock         : in  std_logic                     := 'X';             -- clk
			fir_in_data   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			fir_in_ready  : out std_logic;                                        -- ready
			fir_in_valid  : in  std_logic                     := 'X';             -- valid
			fir_out_data  : out std_logic_vector(31 downto 0);                    -- data
			fir_out_ready : in  std_logic                     := 'X';             -- ready
			fir_out_valid : out std_logic;                                        -- valid
			resetn        : in  std_logic                     := 'X';             -- reset_n
			done          : out std_logic;                                        -- valid
			stall         : in  std_logic                     := 'X'              -- stall
		);
	end component embedded_computer_system_filter_0;

	component embedded_computer_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component embedded_computer_system_jtag_uart;

	component embedded_computer_system_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component embedded_computer_system_onchip_ram;

	component embedded_computer_system_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component embedded_computer_system_pll;

	component embedded_computer_system_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component embedded_computer_system_sdram_controller;

	component embedded_computer_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component embedded_computer_system_sysid_qsys_0;

	component embedded_computer_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                  : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                 : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			buffer_0_avs_cra_address                              : out std_logic_vector(2 downto 0);                     -- address
			buffer_0_avs_cra_write                                : out std_logic;                                        -- write
			buffer_0_avs_cra_read                                 : out std_logic;                                        -- read
			buffer_0_avs_cra_readdata                             : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			buffer_0_avs_cra_writedata                            : out std_logic_vector(63 downto 0);                    -- writedata
			buffer_0_avs_cra_byteenable                           : out std_logic_vector(7 downto 0);                     -- byteenable
			buffer_0_avs_sample_buffer_address                    : out std_logic_vector(8 downto 0);                     -- address
			buffer_0_avs_sample_buffer_write                      : out std_logic;                                        -- write
			buffer_0_avs_sample_buffer_read                       : out std_logic;                                        -- read
			buffer_0_avs_sample_buffer_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			buffer_0_avs_sample_buffer_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			buffer_0_avs_sample_buffer_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			buffer_1_avs_result_buffer_address                    : out std_logic_vector(8 downto 0);                     -- address
			buffer_1_avs_result_buffer_write                      : out std_logic;                                        -- write
			buffer_1_avs_result_buffer_read                       : out std_logic;                                        -- read
			buffer_1_avs_result_buffer_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			buffer_1_avs_result_buffer_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			buffer_1_avs_result_buffer_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                             : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                              : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			onchip_ram_s1_address                                 : out std_logic_vector(11 downto 0);                    -- address
			onchip_ram_s1_write                                   : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                   : out std_logic;                                        -- clken
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_controller_s1_address                           : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                             : out std_logic;                                        -- write
			sdram_controller_s1_read                              : out std_logic;                                        -- read
			sdram_controller_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                        : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_HW_IP_0_avalon_slave_0_address                  : out std_logic_vector(1 downto 0);                     -- address
			TIMER_HW_IP_0_avalon_slave_0_write                    : out std_logic;                                        -- write
			TIMER_HW_IP_0_avalon_slave_0_read                     : out std_logic;                                        -- read
			TIMER_HW_IP_0_avalon_slave_0_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_HW_IP_0_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			TIMER_HW_IP_0_avalon_slave_0_chipselect               : out std_logic;                                        -- chipselect
			VGA_IP_0_avalon_slave_0_address                       : out std_logic_vector(16 downto 0);                    -- address
			VGA_IP_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			VGA_IP_0_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_IP_0_avalon_slave_0_chipselect                    : out std_logic                                         -- chipselect
		);
	end component embedded_computer_system_mm_interconnect_0;

	component embedded_computer_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component embedded_computer_system_irq_mapper;

	component embedded_computer_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component embedded_computer_system_rst_controller;

	component embedded_computer_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component embedded_computer_system_rst_controller_001;

	component embedded_computer_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component embedded_computer_system_rst_controller_002;

	signal filter_0_fir_out_valid                                              : std_logic;                     -- filter_0:fir_out_valid -> buffer_1:result_in_valid
	signal filter_0_fir_out_data                                               : std_logic_vector(31 downto 0); -- filter_0:fir_out_data -> buffer_1:result_in_data
	signal filter_0_fir_out_ready                                              : std_logic;                     -- buffer_1:result_in_ready -> filter_0:fir_out_ready
	signal buffer_0_sample_out_valid                                           : std_logic;                     -- buffer_0:sample_out_valid -> filter_0:fir_in_valid
	signal buffer_0_sample_out_data                                            : std_logic_vector(15 downto 0); -- buffer_0:sample_out_data -> filter_0:fir_in_data
	signal buffer_0_sample_out_ready                                           : std_logic;                     -- filter_0:fir_in_ready -> buffer_0:sample_out_ready
	signal pll_c0_clk                                                          : std_logic;                     -- pll:c0 -> [TIMER_HW_IP_0:clk, VGA_IP_0:CLOCK_controller_50, buffer_0:clock, buffer_1:clock, cpu:clk, filter_0:clock, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_c0_clk, onchip_ram:clk, rst_controller:clk, rst_controller_001:clk, sdram_controller:clk, sysid_qsys_0:clock]
	signal cpu_data_master_readdata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                         : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                         : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                             : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                          : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                               : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                           : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                      : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                         : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata              : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest           : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                  : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                 : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect           : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata             : std_logic_vector(31 downto 0); -- TIMER_HW_IP_0:dout -> mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_readdata
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_address -> TIMER_HW_IP_0:addr
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read                 : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_read -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write                : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_write -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_writedata -> TIMER_HW_IP_0:din
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect                : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_address                   : std_logic_vector(16 downto 0); -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_address -> VGA_IP_0:address_controller_in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_write                     : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_write -> VGA_IP_0:wren_controller
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_writedata -> VGA_IP_0:data_controller_in
	signal mm_interconnect_0_buffer_0_avs_cra_readdata                         : std_logic_vector(63 downto 0); -- buffer_0:avs_cra_readdata -> mm_interconnect_0:buffer_0_avs_cra_readdata
	signal mm_interconnect_0_buffer_0_avs_cra_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:buffer_0_avs_cra_address -> buffer_0:avs_cra_address
	signal mm_interconnect_0_buffer_0_avs_cra_read                             : std_logic;                     -- mm_interconnect_0:buffer_0_avs_cra_read -> buffer_0:avs_cra_read
	signal mm_interconnect_0_buffer_0_avs_cra_byteenable                       : std_logic_vector(7 downto 0);  -- mm_interconnect_0:buffer_0_avs_cra_byteenable -> buffer_0:avs_cra_byteenable
	signal mm_interconnect_0_buffer_0_avs_cra_write                            : std_logic;                     -- mm_interconnect_0:buffer_0_avs_cra_write -> buffer_0:avs_cra_write
	signal mm_interconnect_0_buffer_0_avs_cra_writedata                        : std_logic_vector(63 downto 0); -- mm_interconnect_0:buffer_0_avs_cra_writedata -> buffer_0:avs_cra_writedata
	signal mm_interconnect_0_buffer_1_avs_result_buffer_readdata               : std_logic_vector(31 downto 0); -- buffer_1:avs_result_buffer_readdata -> mm_interconnect_0:buffer_1_avs_result_buffer_readdata
	signal mm_interconnect_0_buffer_1_avs_result_buffer_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:buffer_1_avs_result_buffer_address -> buffer_1:avs_result_buffer_address
	signal mm_interconnect_0_buffer_1_avs_result_buffer_read                   : std_logic;                     -- mm_interconnect_0:buffer_1_avs_result_buffer_read -> buffer_1:avs_result_buffer_read
	signal mm_interconnect_0_buffer_1_avs_result_buffer_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:buffer_1_avs_result_buffer_byteenable -> buffer_1:avs_result_buffer_byteenable
	signal mm_interconnect_0_buffer_1_avs_result_buffer_write                  : std_logic;                     -- mm_interconnect_0:buffer_1_avs_result_buffer_write -> buffer_1:avs_result_buffer_write
	signal mm_interconnect_0_buffer_1_avs_result_buffer_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:buffer_1_avs_result_buffer_writedata -> buffer_1:avs_result_buffer_writedata
	signal mm_interconnect_0_buffer_0_avs_sample_buffer_readdata               : std_logic_vector(31 downto 0); -- buffer_0:avs_sample_buffer_readdata -> mm_interconnect_0:buffer_0_avs_sample_buffer_readdata
	signal mm_interconnect_0_buffer_0_avs_sample_buffer_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:buffer_0_avs_sample_buffer_address -> buffer_0:avs_sample_buffer_address
	signal mm_interconnect_0_buffer_0_avs_sample_buffer_read                   : std_logic;                     -- mm_interconnect_0:buffer_0_avs_sample_buffer_read -> buffer_0:avs_sample_buffer_read
	signal mm_interconnect_0_buffer_0_avs_sample_buffer_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:buffer_0_avs_sample_buffer_byteenable -> buffer_0:avs_sample_buffer_byteenable
	signal mm_interconnect_0_buffer_0_avs_sample_buffer_write                  : std_logic;                     -- mm_interconnect_0:buffer_0_avs_sample_buffer_write -> buffer_0:avs_sample_buffer_write
	signal mm_interconnect_0_buffer_0_avs_sample_buffer_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:buffer_0_avs_sample_buffer_writedata -> buffer_0:avs_sample_buffer_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata               : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                      : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                   : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                          : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                         : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                            : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                                : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                               : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                            : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                             : std_logic_vector(11 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                               : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                               : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_sdram_controller_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                      : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest                   : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                       : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                          : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid                 : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                         : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- buffer_0:done_irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [onchip_ram:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                       : std_logic;                     -- cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_001_reset_out_reset_req                              : std_logic;                     -- rst_controller_001:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_002_reset_out_reset                                  : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv        : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect:inv -> TIMER_HW_IP_0:cs_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv       : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read:inv -> TIMER_HW_IP_0:read_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv      : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write:inv -> TIMER_HW_IP_0:write_n
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv      : std_logic;                     -- mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect:inv -> VGA_IP_0:cs_n
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv                : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv          : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [TIMER_HW_IP_0:reset_n, VGA_IP_0:reset_controller, jtag_uart:rst_n, sdram_controller:reset_n, sysid_qsys_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [buffer_0:resetn, buffer_1:resetn, cpu:reset_n, filter_0:resetn]

begin

	timer_hw_ip_0 : component TIMER_HW_IP
		port map (
			reset_n => rst_controller_reset_out_reset_ports_inv,                            --          reset.reset_n
			clk     => pll_c0_clk,                                                          --          clock.clk
			cs_n    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			addr    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address,              --               .address
			write_n => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv,      --               .write_n
			read_n  => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv,       --               .read_n
			din     => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata,            --               .writedata
			dout    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata              --               .readdata
		);

	vga_ip_0 : component VGA_IP
		port map (
			data_controller_in    => mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata,            -- avalon_slave_0.writedata
			wren_controller       => mm_interconnect_0_vga_ip_0_avalon_slave_0_write,                --               .write
			cs_n                  => mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv, --               .chipselect_n
			address_controller_in => mm_interconnect_0_vga_ip_0_avalon_slave_0_address,              --               .address
			reset_controller      => rst_controller_reset_out_reset_ports_inv,                       --          reset.reset_n
			CLOCK_controller_50   => pll_c0_clk,                                                     --          clock.clk
			VGA_controller_B      => vga_ip_0_conduit_end_vga_b,                                     --    conduit_end.vga_b
			VGA_controller_G      => vga_ip_0_conduit_end_vga_g,                                     --               .vga_g
			VGA_controller_R      => vga_ip_0_conduit_end_vga_r,                                     --               .vga_r
			VGA_controller_VS     => vga_ip_0_conduit_end_vga_vs,                                    --               .vga_vs
			VGA_controller_HS     => vga_ip_0_conduit_end_vga_hs                                     --               .vga_hs
		);

	buffer_0 : component embedded_computer_system_buffer_0
		port map (
			avs_cra_read                 => mm_interconnect_0_buffer_0_avs_cra_read,                 --           avs_cra.read
			avs_cra_write                => mm_interconnect_0_buffer_0_avs_cra_write,                --                  .write
			avs_cra_address              => mm_interconnect_0_buffer_0_avs_cra_address,              --                  .address
			avs_cra_writedata            => mm_interconnect_0_buffer_0_avs_cra_writedata,            --                  .writedata
			avs_cra_byteenable           => mm_interconnect_0_buffer_0_avs_cra_byteenable,           --                  .byteenable
			avs_cra_readdata             => mm_interconnect_0_buffer_0_avs_cra_readdata,             --                  .readdata
			avs_sample_buffer_read       => mm_interconnect_0_buffer_0_avs_sample_buffer_read,       -- avs_sample_buffer.read
			avs_sample_buffer_write      => mm_interconnect_0_buffer_0_avs_sample_buffer_write,      --                  .write
			avs_sample_buffer_address    => mm_interconnect_0_buffer_0_avs_sample_buffer_address,    --                  .address
			avs_sample_buffer_writedata  => mm_interconnect_0_buffer_0_avs_sample_buffer_writedata,  --                  .writedata
			avs_sample_buffer_byteenable => mm_interconnect_0_buffer_0_avs_sample_buffer_byteenable, --                  .byteenable
			avs_sample_buffer_readdata   => mm_interconnect_0_buffer_0_avs_sample_buffer_readdata,   --                  .readdata
			clock                        => pll_c0_clk,                                              --             clock.clk
			done_irq                     => irq_mapper_receiver1_irq,                                --               irq.irq
			resetn                       => rst_controller_001_reset_out_reset_ports_inv,            --             reset.reset_n
			sample_out_data              => buffer_0_sample_out_data,                                --        sample_out.data
			sample_out_ready             => buffer_0_sample_out_ready,                               --                  .ready
			sample_out_valid             => buffer_0_sample_out_valid                                --                  .valid
		);

	buffer_1 : component embedded_computer_system_buffer_1
		port map (
			avs_result_buffer_read       => mm_interconnect_0_buffer_1_avs_result_buffer_read,       -- avs_result_buffer.read
			avs_result_buffer_write      => mm_interconnect_0_buffer_1_avs_result_buffer_write,      --                  .write
			avs_result_buffer_address    => mm_interconnect_0_buffer_1_avs_result_buffer_address,    --                  .address
			avs_result_buffer_writedata  => mm_interconnect_0_buffer_1_avs_result_buffer_writedata,  --                  .writedata
			avs_result_buffer_byteenable => mm_interconnect_0_buffer_1_avs_result_buffer_byteenable, --                  .byteenable
			avs_result_buffer_readdata   => mm_interconnect_0_buffer_1_avs_result_buffer_readdata,   --                  .readdata
			start                        => buffer_1_call_valid,                                     --              call.valid
			busy                         => buffer_1_call_stall,                                     --                  .stall
			clock                        => pll_c0_clk,                                              --             clock.clk
			resetn                       => rst_controller_001_reset_out_reset_ports_inv,            --             reset.reset_n
			result_in_data               => filter_0_fir_out_data,                                   --         result_in.data
			result_in_ready              => filter_0_fir_out_ready,                                  --                  .ready
			result_in_valid              => filter_0_fir_out_valid,                                  --                  .valid
			done                         => buffer_1_return_valid,                                   --            return.valid
			stall                        => buffer_1_return_stall                                    --                  .stall
		);

	cpu : component embedded_computer_system_cpu
		port map (
			clk                                 => pll_c0_clk,                                        --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	filter_0 : component embedded_computer_system_filter_0
		port map (
			start         => filter_0_call_valid,                          --    call.valid
			busy          => filter_0_call_stall,                          --        .stall
			clock         => pll_c0_clk,                                   --   clock.clk
			fir_in_data   => buffer_0_sample_out_data,                     --  fir_in.data
			fir_in_ready  => buffer_0_sample_out_ready,                    --        .ready
			fir_in_valid  => buffer_0_sample_out_valid,                    --        .valid
			fir_out_data  => filter_0_fir_out_data,                        -- fir_out.data
			fir_out_ready => filter_0_fir_out_ready,                       --        .ready
			fir_out_valid => filter_0_fir_out_valid,                       --        .valid
			resetn        => rst_controller_001_reset_out_reset_ports_inv, --   reset.reset_n
			done          => filter_0_return_valid,                        --  return.valid
			stall         => filter_0_return_stall                         --        .stall
		);

	jtag_uart : component embedded_computer_system_jtag_uart
		port map (
			clk            => pll_c0_clk,                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	onchip_ram : component embedded_computer_system_onchip_ram
		port map (
			clk        => pll_c0_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pll : component embedded_computer_system_pll
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_002_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => pll_c1_clk,                                --                    c1.clk
			c2                 => open,                                      --                    c2.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	sdram_controller : component embedded_computer_system_sdram_controller
		port map (
			clk            => pll_c0_clk,                                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_addr,                                      --  wire.export
			zs_ba          => sdram_controller_ba,                                        --      .export
			zs_cas_n       => sdram_controller_cas_n,                                     --      .export
			zs_cke         => sdram_controller_cke,                                       --      .export
			zs_cs_n        => sdram_controller_cs_n,                                      --      .export
			zs_dq          => sdram_controller_dq,                                        --      .export
			zs_dqm         => sdram_controller_dqm,                                       --      .export
			zs_ras_n       => sdram_controller_ras_n,                                     --      .export
			zs_we_n        => sdram_controller_we_n                                       --      .export
		);

	sysid_qsys_0 : component embedded_computer_system_sysid_qsys_0
		port map (
			clock    => pll_c0_clk,                                              --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component embedded_computer_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                         => clk_clk,                                                   --                                       clk_0_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                                --                                          pll_c0.clk
			cpu_reset_reset_bridge_in_reset_reset                 => rst_controller_001_reset_out_reset,                        --                 cpu_reset_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset           => rst_controller_reset_out_reset,                            --           jtag_uart_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                        -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                               => cpu_data_master_address,                                   --                                 cpu_data_master.address
			cpu_data_master_waitrequest                           => cpu_data_master_waitrequest,                               --                                                .waitrequest
			cpu_data_master_byteenable                            => cpu_data_master_byteenable,                                --                                                .byteenable
			cpu_data_master_read                                  => cpu_data_master_read,                                      --                                                .read
			cpu_data_master_readdata                              => cpu_data_master_readdata,                                  --                                                .readdata
			cpu_data_master_write                                 => cpu_data_master_write,                                     --                                                .write
			cpu_data_master_writedata                             => cpu_data_master_writedata,                                 --                                                .writedata
			cpu_data_master_debugaccess                           => cpu_data_master_debugaccess,                               --                                                .debugaccess
			cpu_instruction_master_address                        => cpu_instruction_master_address,                            --                          cpu_instruction_master.address
			cpu_instruction_master_waitrequest                    => cpu_instruction_master_waitrequest,                        --                                                .waitrequest
			cpu_instruction_master_read                           => cpu_instruction_master_read,                               --                                                .read
			cpu_instruction_master_readdata                       => cpu_instruction_master_readdata,                           --                                                .readdata
			buffer_0_avs_cra_address                              => mm_interconnect_0_buffer_0_avs_cra_address,                --                                buffer_0_avs_cra.address
			buffer_0_avs_cra_write                                => mm_interconnect_0_buffer_0_avs_cra_write,                  --                                                .write
			buffer_0_avs_cra_read                                 => mm_interconnect_0_buffer_0_avs_cra_read,                   --                                                .read
			buffer_0_avs_cra_readdata                             => mm_interconnect_0_buffer_0_avs_cra_readdata,               --                                                .readdata
			buffer_0_avs_cra_writedata                            => mm_interconnect_0_buffer_0_avs_cra_writedata,              --                                                .writedata
			buffer_0_avs_cra_byteenable                           => mm_interconnect_0_buffer_0_avs_cra_byteenable,             --                                                .byteenable
			buffer_0_avs_sample_buffer_address                    => mm_interconnect_0_buffer_0_avs_sample_buffer_address,      --                      buffer_0_avs_sample_buffer.address
			buffer_0_avs_sample_buffer_write                      => mm_interconnect_0_buffer_0_avs_sample_buffer_write,        --                                                .write
			buffer_0_avs_sample_buffer_read                       => mm_interconnect_0_buffer_0_avs_sample_buffer_read,         --                                                .read
			buffer_0_avs_sample_buffer_readdata                   => mm_interconnect_0_buffer_0_avs_sample_buffer_readdata,     --                                                .readdata
			buffer_0_avs_sample_buffer_writedata                  => mm_interconnect_0_buffer_0_avs_sample_buffer_writedata,    --                                                .writedata
			buffer_0_avs_sample_buffer_byteenable                 => mm_interconnect_0_buffer_0_avs_sample_buffer_byteenable,   --                                                .byteenable
			buffer_1_avs_result_buffer_address                    => mm_interconnect_0_buffer_1_avs_result_buffer_address,      --                      buffer_1_avs_result_buffer.address
			buffer_1_avs_result_buffer_write                      => mm_interconnect_0_buffer_1_avs_result_buffer_write,        --                                                .write
			buffer_1_avs_result_buffer_read                       => mm_interconnect_0_buffer_1_avs_result_buffer_read,         --                                                .read
			buffer_1_avs_result_buffer_readdata                   => mm_interconnect_0_buffer_1_avs_result_buffer_readdata,     --                                                .readdata
			buffer_1_avs_result_buffer_writedata                  => mm_interconnect_0_buffer_1_avs_result_buffer_writedata,    --                                                .writedata
			buffer_1_avs_result_buffer_byteenable                 => mm_interconnect_0_buffer_1_avs_result_buffer_byteenable,   --                                                .byteenable
			cpu_debug_mem_slave_address                           => mm_interconnect_0_cpu_debug_mem_slave_address,             --                             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                             => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                                .write
			cpu_debug_mem_slave_read                              => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                                .read
			cpu_debug_mem_slave_readdata                          => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                                .readdata
			cpu_debug_mem_slave_writedata                         => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                                .writedata
			cpu_debug_mem_slave_byteenable                        => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                                .byteenable
			cpu_debug_mem_slave_waitrequest                       => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                                .waitrequest
			cpu_debug_mem_slave_debugaccess                       => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                                .debugaccess
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                .chipselect
			onchip_ram_s1_address                                 => mm_interconnect_0_onchip_ram_s1_address,                   --                                   onchip_ram_s1.address
			onchip_ram_s1_write                                   => mm_interconnect_0_onchip_ram_s1_write,                     --                                                .write
			onchip_ram_s1_readdata                                => mm_interconnect_0_onchip_ram_s1_readdata,                  --                                                .readdata
			onchip_ram_s1_writedata                               => mm_interconnect_0_onchip_ram_s1_writedata,                 --                                                .writedata
			onchip_ram_s1_byteenable                              => mm_interconnect_0_onchip_ram_s1_byteenable,                --                                                .byteenable
			onchip_ram_s1_chipselect                              => mm_interconnect_0_onchip_ram_s1_chipselect,                --                                                .chipselect
			onchip_ram_s1_clken                                   => mm_interconnect_0_onchip_ram_s1_clken,                     --                                                .clken
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,                   --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,                     --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                      --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,                  --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,                 --                                                .writedata
			sdram_controller_s1_address                           => mm_interconnect_0_sdram_controller_s1_address,             --                             sdram_controller_s1.address
			sdram_controller_s1_write                             => mm_interconnect_0_sdram_controller_s1_write,               --                                                .write
			sdram_controller_s1_read                              => mm_interconnect_0_sdram_controller_s1_read,                --                                                .read
			sdram_controller_s1_readdata                          => mm_interconnect_0_sdram_controller_s1_readdata,            --                                                .readdata
			sdram_controller_s1_writedata                         => mm_interconnect_0_sdram_controller_s1_writedata,           --                                                .writedata
			sdram_controller_s1_byteenable                        => mm_interconnect_0_sdram_controller_s1_byteenable,          --                                                .byteenable
			sdram_controller_s1_readdatavalid                     => mm_interconnect_0_sdram_controller_s1_readdatavalid,       --                                                .readdatavalid
			sdram_controller_s1_waitrequest                       => mm_interconnect_0_sdram_controller_s1_waitrequest,         --                                                .waitrequest
			sdram_controller_s1_chipselect                        => mm_interconnect_0_sdram_controller_s1_chipselect,          --                                                .chipselect
			sysid_qsys_0_control_slave_address                    => mm_interconnect_0_sysid_qsys_0_control_slave_address,      --                      sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                   => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,     --                                                .readdata
			TIMER_HW_IP_0_avalon_slave_0_address                  => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address,    --                    TIMER_HW_IP_0_avalon_slave_0.address
			TIMER_HW_IP_0_avalon_slave_0_write                    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write,      --                                                .write
			TIMER_HW_IP_0_avalon_slave_0_read                     => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read,       --                                                .read
			TIMER_HW_IP_0_avalon_slave_0_readdata                 => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata,   --                                                .readdata
			TIMER_HW_IP_0_avalon_slave_0_writedata                => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata,  --                                                .writedata
			TIMER_HW_IP_0_avalon_slave_0_chipselect               => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect, --                                                .chipselect
			VGA_IP_0_avalon_slave_0_address                       => mm_interconnect_0_vga_ip_0_avalon_slave_0_address,         --                         VGA_IP_0_avalon_slave_0.address
			VGA_IP_0_avalon_slave_0_write                         => mm_interconnect_0_vga_ip_0_avalon_slave_0_write,           --                                                .write
			VGA_IP_0_avalon_slave_0_writedata                     => mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata,       --                                                .writedata
			VGA_IP_0_avalon_slave_0_chipselect                    => mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect       --                                                .chipselect
		);

	irq_mapper : component embedded_computer_system_irq_mapper
		port map (
			clk           => pll_c0_clk,                         --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	rst_controller : component embedded_computer_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component embedded_computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => pll_c0_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component embedded_computer_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write;

	mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of embedded_computer_system
