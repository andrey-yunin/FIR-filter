-- embedded_computer_system_buffer_0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity embedded_computer_system_buffer_0 is
	port (
		avs_cra_read                 : in  std_logic                     := '0';             --           avs_cra.read
		avs_cra_write                : in  std_logic                     := '0';             --                  .write
		avs_cra_address              : in  std_logic_vector(2 downto 0)  := (others => '0'); --                  .address
		avs_cra_writedata            : in  std_logic_vector(63 downto 0) := (others => '0'); --                  .writedata
		avs_cra_byteenable           : in  std_logic_vector(7 downto 0)  := (others => '0'); --                  .byteenable
		avs_cra_readdata             : out std_logic_vector(63 downto 0);                    --                  .readdata
		avs_sample_buffer_read       : in  std_logic                     := '0';             -- avs_sample_buffer.read
		avs_sample_buffer_write      : in  std_logic                     := '0';             --                  .write
		avs_sample_buffer_address    : in  std_logic_vector(8 downto 0)  := (others => '0'); --                  .address
		avs_sample_buffer_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		avs_sample_buffer_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                  .byteenable
		avs_sample_buffer_readdata   : out std_logic_vector(31 downto 0);                    --                  .readdata
		clock                        : in  std_logic                     := '0';             --             clock.clk
		done_irq                     : out std_logic;                                        --               irq.irq
		resetn                       : in  std_logic                     := '0';             --             reset.reset_n
		sample_out_data              : out std_logic_vector(15 downto 0);                    --        sample_out.data
		sample_out_ready             : in  std_logic                     := '0';             --                  .ready
		sample_out_valid             : out std_logic                                         --                  .valid
	);
end entity embedded_computer_system_buffer_0;

architecture rtl of embedded_computer_system_buffer_0 is
	component sample_buffer_internal is
		port (
			clock                        : in  std_logic                     := 'X';             -- clk
			resetn                       : in  std_logic                     := 'X';             -- reset_n
			sample_out_data              : out std_logic_vector(15 downto 0);                    -- data
			sample_out_ready             : in  std_logic                     := 'X';             -- ready
			sample_out_valid             : out std_logic;                                        -- valid
			done_irq                     : out std_logic;                                        -- irq
			avs_cra_read                 : in  std_logic                     := 'X';             -- read
			avs_cra_write                : in  std_logic                     := 'X';             -- write
			avs_cra_address              : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avs_cra_writedata            : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cra_byteenable           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avs_cra_readdata             : out std_logic_vector(63 downto 0);                    -- readdata
			avs_sample_buffer_read       : in  std_logic                     := 'X';             -- read
			avs_sample_buffer_write      : in  std_logic                     := 'X';             -- write
			avs_sample_buffer_address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			avs_sample_buffer_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_sample_buffer_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_sample_buffer_readdata   : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component sample_buffer_internal;

begin

	sample_buffer_internal_inst : component sample_buffer_internal
		port map (
			clock                        => clock,                        --             clock.clk
			resetn                       => resetn,                       --             reset.reset_n
			sample_out_data              => sample_out_data,              --        sample_out.data
			sample_out_ready             => sample_out_ready,             --                  .ready
			sample_out_valid             => sample_out_valid,             --                  .valid
			done_irq                     => done_irq,                     --               irq.irq
			avs_cra_read                 => avs_cra_read,                 --           avs_cra.read
			avs_cra_write                => avs_cra_write,                --                  .write
			avs_cra_address              => avs_cra_address,              --                  .address
			avs_cra_writedata            => avs_cra_writedata,            --                  .writedata
			avs_cra_byteenable           => avs_cra_byteenable,           --                  .byteenable
			avs_cra_readdata             => avs_cra_readdata,             --                  .readdata
			avs_sample_buffer_read       => avs_sample_buffer_read,       -- avs_sample_buffer.read
			avs_sample_buffer_write      => avs_sample_buffer_write,      --                  .write
			avs_sample_buffer_address    => avs_sample_buffer_address,    --                  .address
			avs_sample_buffer_writedata  => avs_sample_buffer_writedata,  --                  .writedata
			avs_sample_buffer_byteenable => avs_sample_buffer_byteenable, --                  .byteenable
			avs_sample_buffer_readdata   => avs_sample_buffer_readdata    --                  .readdata
		);

end architecture rtl; -- of embedded_computer_system_buffer_0
