-- embedded_computer_system_filter_0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity embedded_computer_system_filter_0 is
	port (
		start         : in  std_logic                     := '0';             --    call.valid
		busy          : out std_logic;                                        --        .stall
		clock         : in  std_logic                     := '0';             --   clock.clk
		fir_in_data   : in  std_logic_vector(15 downto 0) := (others => '0'); --  fir_in.data
		fir_in_ready  : out std_logic;                                        --        .ready
		fir_in_valid  : in  std_logic                     := '0';             --        .valid
		fir_out_data  : out std_logic_vector(31 downto 0);                    -- fir_out.data
		fir_out_ready : in  std_logic                     := '0';             --        .ready
		fir_out_valid : out std_logic;                                        --        .valid
		resetn        : in  std_logic                     := '0';             --   reset.reset_n
		done          : out std_logic;                                        --  return.valid
		stall         : in  std_logic                     := '0'              --        .stall
	);
end entity embedded_computer_system_filter_0;

architecture rtl of embedded_computer_system_filter_0 is
	component fir_filter_internal is
		port (
			clock         : in  std_logic                     := 'X';             -- clk
			resetn        : in  std_logic                     := 'X';             -- reset_n
			fir_in_data   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			fir_in_ready  : out std_logic;                                        -- ready
			fir_in_valid  : in  std_logic                     := 'X';             -- valid
			fir_out_data  : out std_logic_vector(31 downto 0);                    -- data
			fir_out_ready : in  std_logic                     := 'X';             -- ready
			fir_out_valid : out std_logic;                                        -- valid
			start         : in  std_logic                     := 'X';             -- valid
			busy          : out std_logic;                                        -- stall
			done          : out std_logic;                                        -- valid
			stall         : in  std_logic                     := 'X'              -- stall
		);
	end component fir_filter_internal;

begin

	fir_filter_internal_inst : component fir_filter_internal
		port map (
			clock         => clock,         --   clock.clk
			resetn        => resetn,        --   reset.reset_n
			fir_in_data   => fir_in_data,   --  fir_in.data
			fir_in_ready  => fir_in_ready,  --        .ready
			fir_in_valid  => fir_in_valid,  --        .valid
			fir_out_data  => fir_out_data,  -- fir_out.data
			fir_out_ready => fir_out_ready, --        .ready
			fir_out_valid => fir_out_valid, --        .valid
			start         => start,         --    call.valid
			busy          => busy,          --        .stall
			done          => done,          --  return.valid
			stall         => stall          --        .stall
		);

end architecture rtl; -- of embedded_computer_system_filter_0
